library verilog;
use verilog.vl_types.all;
entity tb_DDFS_frequency_converter is
end tb_DDFS_frequency_converter;
